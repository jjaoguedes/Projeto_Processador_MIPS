module dsf_OR(
  input a,
  input b,
  output c
);

assign c = a | b;

endmodule