library verilog;
use verilog.vl_types.all;
entity dsf_ALU_vlg_vec_tst is
end dsf_ALU_vlg_vec_tst;
