library verilog;
use verilog.vl_types.all;
entity dsf_somador_completo_vlg_vec_tst is
end dsf_somador_completo_vlg_vec_tst;
