library verilog;
use verilog.vl_types.all;
entity dsf_Mult2to1_vlg_check_tst is
    port(
        \Out\           : in     vl_logic_vector(0 downto 0);
        sampler_rx      : in     vl_logic
    );
end dsf_Mult2to1_vlg_check_tst;
