library verilog;
use verilog.vl_types.all;
entity dsf_Mult4to1_vlg_vec_tst is
end dsf_Mult4to1_vlg_vec_tst;
